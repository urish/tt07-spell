`default_nettype none
//
`timescale 1ns / 1ps

/* This testbench just instantiates the module and makes some convenient wires
   that can be driven / tested by the cocotb test.py.
*/
module tb ();

  // Dump the signals to a VCD file. You can view it with gtkwave.
  initial begin
    $dumpfile("tb.vcd");
    $dumpvars(0, tb);
    #1;
  end

  // Wire up the inputs and outputs:
  reg clk;
  reg rst_n;
  reg ena;
  wire [7:0] ui_in = {sram_miso, i_reg_sel, i_shift_in, i_dump, i_load, i_step, i_run};
  reg [7:0] uio_in;
  wire [7:0] uo_out;
  wire [7:0] uio_out;
  wire [7:0] uio_oe;

  reg i_run;
  reg i_step;
  reg i_load;
  reg i_dump;
  reg i_shift_in;
  reg [1:0] i_reg_sel;

  wire o_cpu_sleep = uo_out[0];
  wire o_cpu_stop = uo_out[1];
  wire o_cpu_wait_delay = uo_out[2];
  wire o_shift_out = uo_out[3];

  reg sram_miso;
  wire sram_cs = uo_out[5];
  wire sram_sclk = uo_out[6];
  wire sram_mosi = uo_out[7];

  // Replace tt_um_example with your module name:
  tt_um_urish_spell user_project (

      // Include power ports for the Gate Level test:
`ifdef GL_TEST
      .VPWR(1'b1),
      .VGND(1'b0),
`endif

      .ui_in  (ui_in),    // Dedicated inputs
      .uo_out (uo_out),   // Dedicated outputs
      .uio_in (uio_in),   // IOs: Input path
      .uio_out(uio_out),  // IOs: Output path
      .uio_oe (uio_oe),   // IOs: Enable path (active high: 0=input, 1=output)
      .ena    (ena),      // enable - goes high when design is selected
      .clk    (clk),      // clock
      .rst_n  (rst_n)     // not reset
  );

endmodule
